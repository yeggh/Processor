constant_2_inst : constant_2 PORT MAP (
		result	 => result_sig
	);
