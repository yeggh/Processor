constant_3_inst : constant_3 PORT MAP (
		result	 => result_sig
	);
