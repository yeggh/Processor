constant_0_4bits_inst : constant_0_4bits PORT MAP (
		result	 => result_sig
	);
