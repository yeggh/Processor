ADD_SUB16bits_inst : ADD_SUB16bits PORT MAP (
		add_sub	 => add_sub_sig,
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		result	 => result_sig
	);
