CMP_wizard_inst : CMP_wizard PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		agb	 => agb_sig,
		alb	 => alb_sig
	);
