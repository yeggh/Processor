const_3_inst : const_3 PORT MAP (
		result	 => result_sig
	);
