opcode_0_wizard_inst : opcode_0_wizard PORT MAP (
		result	 => result_sig
	);
