constant_6_inst : constant_6 PORT MAP (
		result	 => result_sig
	);
