wizard_const_adder_inst : wizard_const_adder PORT MAP (
		datab	 => datab_sig,
		result	 => result_sig
	);
