ADD_SUB_wizard_inst : ADD_SUB_wizard PORT MAP (
		add_sub	 => add_sub_sig,
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		result	 => result_sig
	);
