constant_0_8bits_inst : constant_0_8bits PORT MAP (
		result	 => result_sig
	);
