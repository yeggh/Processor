const_2_inst : const_2 PORT MAP (
		result	 => result_sig
	);
