opcode_sub_inst : opcode_sub PORT MAP (
		dataa	 => dataa_sig,
		result	 => result_sig
	);
