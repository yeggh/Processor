constant_1_16bits_inst : constant_1_16bits PORT MAP (
		result	 => result_sig
	);
