const_6_inst : const_6 PORT MAP (
		result	 => result_sig
	);
