constant_1_32bits_inst : constant_1_32bits PORT MAP (
		result	 => result_sig
	);
