SHIFT_wizard_inst : SHIFT_wizard PORT MAP (
		data	 => data_sig,
		direction	 => direction_sig,
		distance	 => distance_sig,
		result	 => result_sig
	);
