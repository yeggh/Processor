constant_0_32bits_inst : constant_0_32bits PORT MAP (
		result	 => result_sig
	);
