const_1_inst : const_1 PORT MAP (
		result	 => result_sig
	);
